/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_linux (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 732;

    const logic [RomSize-1:0][63:0] mem = {
        64'h000000ff_f0c2c004,
        64'h000000ff_f0c2c003,
        64'h000000ff_f0c2c001,
        64'h000000ff_f0c2c005,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_00292520,
        64'h00000000_00000028,
        64'h20736b63_6f6c6220,
        64'h00000000_20666f20,
        64'h0000206b_636f6c62,
        64'h20676e69_79706f63,
        64'h00000000_00000008,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00746669_68732d67,
        64'h65720073_74707572,
        64'h7265746e_6900746e,
        64'h65726170_2d747075,
        64'h72726574_6e690064,
        64'h65657073_2d746e65,
        64'h72727563_00736567,
        64'h6e617200_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'ha9000000_04000000,
        64'h03000000_01000000,
        64'h1d010000_04000000,
        64'h03000000_07000000,
        64'h0a010000_04000000,
        64'h03000000_00000004,
        64'h00000000_000010f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h09000000_02000000,
        64'h0b000000_02000000,
        64'hec000000_10000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00303030_30303131,
        64'h66666640_63696c70,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'h00010000_08000000,
        64'h03000000_00000c00,
        64'h00000000_000002f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h07000000_02000000,
        64'h03000000_02000000,
        64'hec000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000000_30303030,
        64'h32303166_66664074,
        64'h6e696c63_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_00010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h000000f1_ff000000,
        64'h5b000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_ec000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00303030,
        64'h30303031_66666640,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h00000000_e2000000,
        64'h04000000_03000000,
        64'h01000000_d7000000,
        64'h04000000_03000000,
        64'h01000000_c6000000,
        64'h04000000_03000000,
        64'h00c20100_b8000000,
        64'h04000000_03000000,
        64'h80f0fa02_3f000000,
        64'h04000000_03000000,
        64'h00400d00_00000000,
        64'h00c0c2f0_ff000000,
        64'h5b000000_10000000,
        64'h03000000_00303535,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00303030_63326330,
        64'h66666640_74726175,
        64'h01000000_b1000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h5b000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_4f000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_a9000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_79000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_70000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_66000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h5f000000_05000000,
        64'h03000000_00000000,
        64'h5b000000_04000000,
        64'h03000000_00757063,
        64'h4f000000_04000000,
        64'h03000000_80f0fa02,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'he1f50500_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd4040000_28010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h0c050000_38000000,
        64'h34060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000a0d,
        64'h0a0d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d2020,
        64'h20202020_20202020,
        64'h34202f20_426b2034,
        64'h36202020_3a636f73,
        64'h7341202f_20657a69,
        64'h53202032_4c0a0d20,
        64'h20202020_20202020,
        64'h2034202f_20426b20,
        64'h38202020_203a636f,
        64'h73734120_2f20657a,
        64'h69532035_314c0a0d,
        64'h20202020_20202020,
        64'h20203420_2f20426b,
        64'h20382020_20203a63,
        64'h6f737341_202f2065,
        64'h7a695320_44314c0a,
        64'h0d202020_20202020,
        64'h20202034_202f2042,
        64'h6b203631_2020203a,
        64'h636f7373_41202f20,
        64'h657a6953_2049314c,
        64'h0a0d2020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20200a0d_20202020,
        64'h20202020_20202020,
        64'h20202020_424d2034,
        64'h32303120_20202020,
        64'h20202020_3a657a69,
        64'h53204d41_52440a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202068_73656d5f,
        64'h64322020_20202020,
        64'h20202020_203a6b72,
        64'h6f777465_4e0a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20206e77_6f6e6b6e,
        64'h55202020_20202020,
        64'h20203a71_65724620,
        64'h65726f43_0a0d2020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20312020_20202020,
        64'h20202020_20203a73,
        64'h65726f43_230a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20203120_20202020,
        64'h20202020_203a7365,
        64'h6c69542d_59230a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202031_20202020,
        64'h20202020_20203a73,
        64'h656c6954_2d58230a,
        64'h0d202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h200a0d20_20202020,
        64'h20202020_20202020,
        64'h20202020_20203232,
        64'h3a38313a_31312032,
        64'h32303220_33312072,
        64'h614d2020_20202020,
        64'h20203a65_74614420,
        64'h646c6975_420a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h2020296e_6f697461,
        64'h6c756d69_53282065,
        64'h6e6f4e20_20202020,
        64'h2020203a_6472616f,
        64'h42204147_50460a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h0a0d2020_20202020,
        64'h20202020_20202020,
        64'h20202020_20273133,
        64'h66376437_35302762,
        64'h20202020_3a6e6f69,
        64'h73726556_20656e61,
        64'h6972410a_0d202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h27646166_61343464,
        64'h33276220_3a6e6f69,
        64'h73726556_206e6f74,
        64'h69506e65_704f0a0d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h0a0d2d2d_20202020,
        64'h20206d72_6f667461,
        64'h6c502065_6e616972,
        64'h412b6e6f_7469506e,
        64'h65704f20_20202020,
        64'h2d2d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d0a0d,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h80820141_450160a2,
        64'hcfdff0ef_057e65a1,
        64'h45058e7f_f0efb465,
        64'h05130000_15178f3f,
        64'hf0ef15a5_05130000,
        64'h05178a5f_f0efe406,
        64'h38050513_20058593,
        64'h114101c9_c53765f1,
        64'hb395917f_f0efe2e5,
        64'h05130000_1517bbd9,
        64'hbc850513_00001517,
        64'ha39ff0ef_854a933f,
        64'hf0efc8a5_05130000,
        64'h151793ff_f0efc7e5,
        64'h05130000_1517bbfd,
        64'hbf050513_00001517,
        64'ha61ff0ef_852695bf,
        64'hf0efcb25_05130000,
        64'h1517967f_f0efca65,
        64'h05130000_1517c929,
        64'h84aac9bf_f0ef8552,
        64'h8656020b_2583983f,
        64'hf0efc2a5_05130000,
        64'h151798ff_f0efe8e5,
        64'h05130000_1517f579,
        64'h10e30804_84939a3f,
        64'hf0ef2905_c4c50513,
        64'h00001517_ff999be3,
        64'hb05ff0ef_09850009,
        64'hc5039bff_f0efeae5,
        64'h05130000_1517ad7f,
        64'hf0ef6888_9d1ff0ef,
        64'heb050513_00001517,
        64'hae9ff0ef_64889e3f,
        64'hf0efeb25_05130000,
        64'h1517afbf_f0ef0604,
        64'h8c930184_89936088,
        64'h9fdff0ef_ebc50513,
        64'h00001517_fe999be3,
        64'hb5dff0ef_09850009,
        64'hc503ff04_8993a1bf,
        64'hf0efeba5_05130000,
        64'h1517ff89_99e3b7bf,
        64'hf0ef0985_0007c503,
        64'h013c87b3_4981a3bf,
        64'hf0effe04_8c93ebe5,
        64'h05130000_1517b9bf,
        64'hf0ef0ff9_7513a53f,
        64'hf0efeba5_05130000,
        64'h15174b91_4c411005,
        64'h1e631004_892a8b0a,
        64'hd91ff0ef_850a4605,
        64'h71010489_2583a7bf,
        64'hf0efd225_05130000,
        64'h1517b51f_f0ef4556,
        64'ha8dff0ef_ed450513,
        64'h00001517_b63ff0ef,
        64'h4546a9ff_f0efec65,
        64'h05130000_1517bb7f,
        64'hf0ef6526_ab1ff0ef,
        64'heb850513_00001517,
        64'hbc9ff0ef_7502ac3f,
        64'hf0efeba5_05130000,
        64'h1517bdbf_f0ef6562,
        64'had5ff0ef_eb450513,
        64'h00001517_babff0ef,
        64'h4552ae7f_f0efeb65,
        64'h05130000_1517bbdf,
        64'hf0ef4542_af9ff0ef,
        64'heb850513_00001517,
        64'hbcfff0ef_4532b0bf,
        64'hf0efeba5_05130000,
        64'h1517be1f_f0ef4522,
        64'hb1dff0ef_ebc50513,
        64'h00001517_c35ff0ef,
        64'h6502b2ff_f0efebe5,
        64'h05130000_1517b3bf,
        64'hf0efeaa5_05130000,
        64'h1517bf59_54f9b4bf,
        64'hf0efdf25_05130000,
        64'h1517c63f_f0ef8526,
        64'hb5dff0ef_eb450513,
        64'h00001517_b69ff0ef,
        64'hea850513_00001517,
        64'hc90584aa_890ae9ff,
        64'hf0ef850a_45854605,
        64'h7101b87f_f0efde65,
        64'h05130000_15178082,
        64'h61256ca2_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_64468526,
        64'h60e6fa04_011354fd,
        64'hbb5ff0ef_ecc50513,
        64'h00001517_c905ecff,
        64'hf0ef8aae_8a2a1080,
        64'he466e862_ec5ef05a,
        64'hfc4ee0ca_e4a6ec86,
        64'hf456f852_e8a2711d,
        64'hb7bd2c05_be9ff0ef,
        64'hec850513_00001517,
        64'hb7a10b85_20048493,
        64'hff5799e3_e29007a1,
        64'h00e786b3_621000f4,
        64'h86334781_974e009b,
        64'h97139c29_c19ff0ef,
        64'hf2850513_00001517,
        64'h9c29c79f_f0ef0325,
        64'h553b4585_036a053b,
        64'h9c29c37f_f0eff365,
        64'h05130000_15179c29,
        64'hc97ff0ef_854a9c29,
        64'h4585c4ff_f0eff465,
        64'h05130000_15179c29,
        64'hcafff0ef_855a0005,
        64'h041b4585_c69ff0ef,
        64'hf5050513_00001517,
        64'h09841263_060c1363,
        64'h034b7c3b_80826161,
        64'h45016c02_6ba26b42,
        64'h6ae27a02_79a27942,
        64'h74e26406_60a6c9bf,
        64'hf0eff425_05130000,
        64'h1517032b_6563000b,
        64'h8b1b2000_0a930640,
        64'h0a134401_4b8194ae,
        64'h893289aa_e062e85a,
        64'he486e45e_ec56f052,
        64'hf44ef84a_e0a21592,
        64'h80dd45bd_02059493,
        64'hfc26715d_80820141,
        64'h450160a2_ce9ff0ef,
        64'he406fb45_05131141,
        64'h00001517_8082557d,
        64'hb7d900d7_00230785,
        64'h00f60733_06c82683,
        64'hff698b05_5178b77d,
        64'hd6b80785_00074703,
        64'h00f50733_80824501,
        64'hd3b84719_dbb8577d,
        64'h200007b7_02b6e163,
        64'h0007869b_20000837,
        64'h20000537_fff58b85,
        64'h537c2000_0737d3b8,
        64'h200007b7_10600713,
        64'hfff537fd_00010320,
        64'h079304b7_61630007,
        64'h871b4781_200006b7,
        64'hdbb85779_200007b7,
        64'h06b7ee63_10000793,
        64'h80826105_64a2d3b8,
        64'h4719dbb8_64420ff4,
        64'h7513577d_200007b7,
        64'h60e2d97f_f0ef03e5,
        64'h05130000_1517eaff,
        64'hf0ef9101_15024088,
        64'hdadff0ef_05c50513,
        64'h00001517_e3958b85,
        64'h240153fc_57e0ff65,
        64'h8b050647_849353f8,
        64'hd3b81060_07132000,
        64'h07b7fff5_37fd0001,
        64'h06400793_d7a8dbb8,
        64'h5779e426_e822ec06,
        64'h200007b7_1101bbc5,
        64'h610508a5_05130000,
        64'h151764a2_60e26442,
        64'hd03c4799_e09ff0ef,
        64'h0b050513_00001517,
        64'hf21ff0ef_91010204,
        64'h95132481_e21ff0ef,
        64'h0a850513_00001517,
        64'h5064d03c_16600793,
        64'he35ff0ef_0dc50513,
        64'h00001517_f4dff0ef,
        64'h91010204_95132481,
        64'he4dff0ef_0d450513,
        64'h00001517_5064d03c,
        64'h10400793_20000437,
        64'hfff537fd_000147a9,
        64'hc3b84729_200007b7,
        64'he75ff0ef_e426e822,
        64'hec060f45_05131101,
        64'h00001517_80822501,
        64'h41088082_c10c8082,
        64'h61054509_60e2e1ff,
        64'hf0ef0091_4503e27f,
        64'hf0ef0081_4503ed9f,
        64'hf0efec06_002c1101,
        64'h80826145_45416942,
        64'h64e27402_70a2ff24,
        64'h10e3e4bf_f0ef0091,
        64'h4503e53f_f0ef3461,
        64'h00814503_f07ff0ef,
        64'h0ff57513_002c0084,
        64'hd5335961_03800413,
        64'h84aaf406_e84aec26,
        64'hf0227179_80826145,
        64'h45216942_64e27402,
        64'h70a2ff24_10e3e8ff,
        64'hf0ef0091_4503e97f,
        64'hf0ef3461_00814503,
        64'hf4bff0ef_0ff57513,
        64'h002c0084_d53b5961,
        64'h446184aa_f406e84a,
        64'hec26f022_71798082,
        64'h612169e2_854e6b02,
        64'h6aa26a42_790274a2,
        64'h744270e2_fd5913e3,
        64'h397d85d2_eddff0ef,
        64'h0007c503_97ba8bbd,
        64'h02d7d7bb_29856ce7,
        64'h07130000_071702ba,
        64'h706300d7_f4630364,
        64'h543b0009_0a1b0284,
        64'hf4bb0004_069b0004,
        64'h879b5afd_4b294981,
        64'h4925a004_041384aa,
        64'he852fc06_e05ae456,
        64'hec4ef04a_f4263b9a,
        64'hd437f822_71398082,
        64'h00f58023_0007c783,
        64'h00e580a3_97aa8111,
        64'h00074703_973e00f5,
        64'h77137327_87930000,
        64'h0797b7c5_f5dff0ef,
        64'h853e8082_610564a2,
        64'h644260e2_e791fff7,
        64'hc7830084_87b30405,
        64'h0004051b_440184aa,
        64'hec06e426_e8221101,
        64'h808200e7_80230200,
        64'h071354a7_b7830000,
        64'h179700f7_0023478d,
        64'h00a68023_0ff57513,
        64'h00c78023_0085551b,
        64'h0ff57613_07ba30b7,
        64'h879303ff_c7b700f7,
        64'h0023f800_07930006,
        64'h802357a7_b7030000,
        64'h179757a7_b6830000,
        64'h179702b5_553b0045,
        64'h959b8082_00a78023,
        64'h07ba30b7_879303ff,
        64'hc7b7dbe5_0207f793,
        64'h0007c783_59c7b783,
        64'h00001797_80820205,
        64'h75130007_c5035ae7,
        64'hb7830000_17978082,
        64'h0ff57513_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00048067,
        64'h01f49493_0010049b,
        64'hd6058593_00001597,
        64'hf1402573_ff2496e3,
        64'h00100493_0004a903,
        64'h04048493_01a49493,
        64'h0210049b_0924a4af,
        64'h00190913_04048493,
        64'h01a49493_0210049b,
        64'hff2496e3_f14024f3,
        64'h0004a903_04048493,
        64'h01a49493_0210049b,
        64'h07d000ef_01a11113,
        64'h0210011b_01249863,
        64'hf1402973_00000493
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
